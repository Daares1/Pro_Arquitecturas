--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.Std_Logic_1164.all;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ENTITY Configurable_U11 IS
  PORT(
      I : IN std_logic;
      O : OUT std_logic
  );
END Configurable_U11;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ARCHITECTURE structure OF Configurable_U11 IS
BEGIN
    O <= NOT(I);
END structure;
--------------------------------------------------------------------------------
