--------------------------------------------------------------------------------
-- SubModule MUX
-- Created   22/05/2014 08:27:30 p.m.
--------------------------------------------------------------------------------
Library IEEE;
Use IEEE.Std_Logic_1164.all;

entity MUX is port
   (
     S       : in    std_logic_vector(2 downto 0);
     DH      : in    std_logic;
     DG      : in    std_logic;
     DF      : in    std_logic;
     DE      : in    std_logic;
     DD      : in    std_logic;
     DC      : in    std_logic;
     DB      : in    std_logic;
     DA      : in    std_logic;
     Y       : out   std_logic
   );

end MUX;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
architecture Structure of MUX is

-- Component Declarations

-- Signal Declarations

begin

end Structure;
--------------------------------------------------------------------------------
